module i2o_sequencer (
	input clk,
	input rst,  // Asynchronous reset active low

);

endmodule