module sha256_preprocessor (
  input clk,
  input rst,


);

endmodule